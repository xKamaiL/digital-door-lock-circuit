library verilog;
use verilog.vl_types.all;
entity look_door_01_vlg_check_tst is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        A3              : in     vl_logic;
        A4              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end look_door_01_vlg_check_tst;
