library verilog;
use verilog.vl_types.all;
entity look_door_01_vlg_vec_tst is
end look_door_01_vlg_vec_tst;
